//-------------------------------------------------------------------------
// Module Name: ahb_slave
// The Slave module of AHB Protocol
// Author: WangFW modified by William Inselberger and Leonardo Guedes
//-------------------------------------------------------------------------
// Date: 2020-11-1 and modified on 2024-05
// Basic features about read and write
// Date: 2020-11-1
// New features: wait state, burst
//-------------------------------------------------------------------------

module ahbslave(
  input hclk,
  input hresetn,
  input hsel,
  input [9:0] haddr,
  input hwrite,
  input [2:0] hsize,
  input [2:0] hburst,
  input [3:0] hprot,
  input [1:0] htrans,
  input hmastlock,
  input hready,
  input [7:0] hwdata,
  input [9:0]displaysel,
  output reg hreadyout,
  output reg hresp,
  output reg [7:0] hrdata,
  output [7:0] memo

);

//----------------------------------------------------------------------
// The definitions for intern registers for data storge
//----------------------------------------------------------------------
reg [7:0] mem [2**10-1:0];
reg [9:0] waddr;
reg [9:0] raddr;

//----------------------------------------------------------------------
// The definition for state machine
//----------------------------------------------------------------------
reg [1:0] state;
reg [1:0] next_state;
localparam idle = 2'b00,s1 = 2'b01,WRITE = 2'b10,READ = 2'b11;


assign estadoslave=state;
//----------------------------------------------------------------------
// The definition for burst feature
//----------------------------------------------------------------------
reg single_flag;
reg incr_flag;
reg wrap4_flag;
reg incr4_flag;
reg wrap8_flag;
reg incr8_flag;
reg wrap16_flag;
reg incr16_flag;
assign memo=mem[displaysel];
integer i;

//----------------------------------------------------------------------
// The state machine
//----------------------------------------------------------------------
//initial begin
//
//for(i=0;i<=1023;i=i+1) mem[i]=0;
//
//end

always @(posedge hclk, negedge hresetn) begin
  if(!hresetn) begin
		state <= idle;
  end
  else begin
    state <= next_state;
  end
end

always @(*) begin
  case(state)
    idle: begin
      single_flag = 1'b0;
      incr_flag = 1'b0;
      wrap4_flag = 1'b0;
      incr4_flag = 1'b0;
      wrap8_flag = 1'b0;
      incr8_flag = 1'b0;
      wrap16_flag = 1'b0;
      incr16_flag = 1'b0;
      if(hsel == 1'b1) begin
        next_state = s1;
      end
      else begin
        next_state = idle;
      end
    end
    s1: begin
      case(hburst)
        // single transfer burst
        3'b000: begin  
          single_flag = 1'b1;
          incr_flag = 1'b0;
          wrap4_flag = 1'b0;
          incr4_flag = 1'b0;
          wrap8_flag = 1'b0;
          incr8_flag = 1'b0;
          wrap16_flag = 1'b0;
          incr16_flag = 1'b0;
        end
        // incrementing burst of undefined length
        3'b001: begin  
          single_flag = 1'b0;
          incr_flag = 1'b1;
          wrap4_flag = 1'b0;
          incr4_flag = 1'b0;
          wrap8_flag = 1'b0;
          incr8_flag = 1'b0;
          wrap16_flag = 1'b0;
          incr16_flag = 1'b0;
        end
        // 4-beat wrapping burst
        3'b010: begin  
          single_flag = 1'b0;
          incr_flag = 1'b0;
          wrap4_flag = 1'b1;
          incr4_flag = 1'b0;
          wrap8_flag = 1'b0;
          incr8_flag = 1'b0;
          wrap16_flag = 1'b0;
          incr16_flag = 1'b0;
			 
        end
        // 4-beat incrementing burst
        3'b011: begin  
          single_flag = 1'b0;
          incr_flag = 1'b0;
          wrap4_flag = 1'b0;
          incr4_flag = 1'b1;
          wrap8_flag = 1'b0;
          incr8_flag = 1'b0;
          wrap16_flag = 1'b0;
          incr16_flag = 1'b0;
        end
        // 8-beat wrapping burst
        3'b100: begin  
          single_flag = 1'b0;
          incr_flag = 1'b0;
          wrap4_flag = 1'b0;
          incr4_flag = 1'b0;
          wrap8_flag = 1'b1;
          incr8_flag = 1'b0;
          wrap16_flag = 1'b0;
          incr16_flag = 1'b0;
        end
        // 8-beat incrementing burst
        3'b101: begin  
          single_flag = 1'b0;
          incr_flag = 1'b0;
          wrap4_flag = 1'b0;
          incr4_flag = 1'b0;
          wrap8_flag = 1'b0;
          incr8_flag = 1'b1;
          wrap16_flag = 1'b0;
          incr16_flag = 1'b0;
        end
        // 16-beat wrapping burst
        3'b110: begin  
          single_flag = 1'b0;
          incr_flag = 1'b0;
          wrap4_flag = 1'b0;
          incr4_flag = 1'b0;
          wrap8_flag = 1'b0;
          incr8_flag = 1'b0;
          wrap16_flag = 1'b1;
          incr16_flag = 1'b0;
        end
        // 16-beat incrementing burst
        3'b111: begin  
          single_flag = 1'b0;
          incr_flag = 1'b0;
          wrap4_flag = 1'b0;
          incr4_flag = 1'b0;
          wrap8_flag = 1'b0;
          incr8_flag = 1'b0;
          wrap16_flag = 1'b0;
          incr16_flag = 1'b1;
        end
        // default
        default: begin  
          single_flag = 1'b0;
          incr_flag = 1'b0;
          wrap4_flag = 1'b0;
          incr4_flag = 1'b0;
          wrap8_flag = 1'b0;
          incr8_flag = 1'b0;
          wrap16_flag = 1'b0;
          incr16_flag = 1'b0;
        end
      endcase
		
		if(htrans!=01) begin
			if(hwrite == 1'b1) begin
				next_state = WRITE;
			end
			else if(hwrite == 1'b0) begin
				next_state = READ;
			end
			else begin
				next_state = s1;
			end
		end
		else begin
			next_state=state;
		end
    end
    WRITE: begin
      case(hburst)
        // single transfer burst
        3'b000: begin  
          if(hsel == 1'b1) begin
            next_state = s1;
          end
          else begin
            next_state = idle;
          end
        end
        // incrementing burst of undefined length
        3'b001: begin  
          next_state = WRITE;
        end
        // 4-beat wrapping burst
        3'b010: begin  
          next_state = WRITE;
        end
        // 4-beat incrementing burst
        3'b011: begin  
          next_state = WRITE;
        end
        // 8-beat wrapping burst
        3'b100: begin  
          next_state = WRITE;
        end
        // 8-beat incrementing burst
        3'b101: begin  
          next_state = WRITE;
        end
        // 16-beat wrapping burst
        3'b110: begin  
          next_state = WRITE;
        end
        // 16-beat incrementing burst
        3'b111: begin  
          next_state = WRITE;
        end
        // default
        default: begin  
          if(hsel == 1'b1) begin
            next_state = s1;
          end
          else begin
            next_state = idle;
          end
        end
      endcase
    end
    READ: begin
      case(hburst)
        // single transfer burst
        3'b000: begin  
          if(hsel == 1'b1) begin
            next_state = s1;
          end
          else begin
            next_state = idle;
          end
        end
        // incrementing burst of undefined length
        3'b001: begin  
          next_state = READ;
        end
        // 4-beat wrapping burst
        3'b010: begin  
          next_state = READ;
        end
        // 4-beat incrementing burst
        3'b011: begin  
          next_state = READ;
        end
        // 8-beat wrapping burst
        3'b100: begin  
          next_state = READ;
        end
        // 8-beat incrementing burst
        3'b101: begin  
          next_state = READ;
        end
        // 16-beat wrapping burst
        3'b110: begin  
          next_state = READ;
        end
        // 16-beat incrementing burst
        3'b111: begin  
          next_state = READ;
        end
        // default
        default: begin  
          if(hsel == 1'b1) begin
            next_state = s1;
          end
          else begin
            next_state = idle;
          end
        end
      endcase
    end
    default: begin
      next_state = idle;
    end
  endcase
end

always @(posedge hclk, negedge hresetn) begin
  if(!hresetn) begin
    hreadyout <= 1'b0;
    hresp <= 1'b0;
    hrdata <= 8'h0_0;
    waddr <= 10'b00_0000_0000;
    raddr <= 10'b00_0000_0000;
	 //for(i=0;i<=1023;i=i+1) mem[i]=0;
  end
  else begin
    case(next_state)
      idle: begin
        hreadyout <= 1'b0;
        hresp <= 1'b0;
        hrdata <= hrdata;
        waddr <= waddr;
        raddr <= raddr;
		  

      end
      s1: begin
        hreadyout <= 1'b0;
        hresp <= 1'b0;
        hrdata <= hrdata;
        waddr <= haddr;
        raddr <= haddr;
		

      end
      WRITE: begin
        case({single_flag,incr_flag,wrap4_flag,incr4_flag,wrap8_flag,incr8_flag,wrap16_flag,incr16_flag})
          // single transfer
          8'b1000_0000: begin
            hreadyout <= 1'b1;
            hresp <= 1'b0;
            mem[waddr] <= hwdata;
          end
          // incre
          8'b0100_0000: begin
            hreadyout <= 1'b1;
            hresp <= 1'b0;
            mem[waddr] <= hwdata;
            waddr <= waddr + 1'b1;
          end
          // wrap 4
          8'b0010_0000: begin

            hresp <= 1'b0;

            if(waddr < haddr+3) begin
              mem[waddr] <= hwdata;
              waddr <= waddr + 1'b1;
				  hreadyout <= 1'b0;
	
				 
            end
            else begin
				/*mem[waddr] <= hwdata;
              waddr <= haddr;*/
				  hreadyout <= 1'b1;
				 
            end
          end
          // incre 4
          8'b0001_0000: begin
           
            hresp <= 1'b0;
				if(waddr>hwdata + 2) hreadyout<=1;
				else  hreadyout <= 1'b0;
            mem[waddr] <= hwdata;
            waddr <= waddr + 1'b1;
				
          end
          // wrap 8
          8'b0000_1000: begin
            hreadyout <= 1'b1;
            hresp <= 1'b0;
            if(waddr < (haddr + 3'd7)) begin
              mem[waddr] <= hwdata;
              waddr <= waddr + 1'b1;
            end
            else begin
              mem[waddr] <= hwdata;
              waddr <= haddr;
            end
          end
          // incre 8
          8'b0000_0100: begin
            hreadyout <= 1'b1;
            hresp <= 1'b0;
            mem[waddr] <= hwdata;
            waddr <= waddr + 1'b1;
          end
          // wrap 16
          8'b0000_0010: begin
            hreadyout <= 1'b1;
            hresp <= 1'b0;
            if(waddr < (haddr + 4'd15)) begin
              mem[waddr] <= hwdata;
              waddr <= waddr + 1'b1;
            end
            else begin
              mem[waddr] <= hwdata;
              waddr <= haddr;
            end
          end
          // incre 16
          8'b0000_0001: begin
            hreadyout <= 1'b1;
            hresp <= 1'b0;
            mem[waddr] <= hwdata;
            waddr <= waddr + 1'b1;
          end
          // default
          default: begin
            hreadyout <= 1'b1;
            hresp <= 1'b0;
          end
        endcase
      end
      READ: begin
        case({single_flag,incr_flag,wrap4_flag,incr4_flag,wrap8_flag,incr8_flag,wrap16_flag,incr16_flag})
          // single transfer
          8'b1000_0000: begin
            hreadyout <= 1'b1;
            hresp <= 1'b0;
            hrdata <= mem[raddr];
          end
          // incre
          8'b0100_0000: begin
            hreadyout <= 1'b1;
            hresp <= 1'b0;
            hrdata <= mem[raddr];
            raddr <= raddr + 1'b1;
          end
          // wrap 4
          8'b0010_0000: begin
          
            hresp <= 1'b0;
            if(raddr < (haddr + 2'd3)) begin
              hrdata <= mem[raddr];
              raddr <= raddr + 1'b1;
				  hreadyout <= 1'b0;
            end
            else begin
             // hrdata <= mem[raddr];
             // raddr <= haddr;
				 hreadyout <= 1'b1;
            end
          end
          // incre 4
          8'b0001_0000: begin
            hreadyout <= 1'b1;
            hresp <= 1'b0;
            hrdata <= mem[raddr];
            raddr <= raddr + 1'b1;
          end
          // wrap 8
          8'b0000_1000: begin
            hreadyout <= 1'b1;
            hresp <= 1'b0;
            if(raddr < (haddr + 3'd7)) begin
              hrdata <= mem[raddr];
              raddr <= raddr + 1'b1;
            end
            else begin
              hrdata <= mem[raddr];
              raddr <= haddr;
            end
          end
          // incre 8
          8'b0000_0100: begin
            hreadyout <= 1'b1;
            hresp <= 1'b0;
            hrdata <= mem[raddr];
            raddr <= raddr + 1'b1;
          end
          // wrap 16
          8'b0000_0010: begin
            hreadyout <= 1'b1;
            hresp <= 1'b0;
            if(raddr < (haddr + 4'd15)) begin
              hrdata <= mem[raddr];
              raddr <= raddr + 1'b1;
            end
            else begin
              hrdata <= mem[raddr];
              raddr <= haddr;
            end
          end
          // incre 16
          8'b0000_0001: begin
            hreadyout <= 1'b1;
            hresp <= 1'b0;
            hrdata <= mem[raddr];
            raddr <= raddr + 1'b1;
          end
          // default
          default: begin
            hreadyout <= 1'b1;
            hresp <= 1'b0;
          end
        endcase
      end
      default: begin
        hreadyout <= 1'b0;
        hresp <= 1'b0;
        hrdata <= hrdata;
        waddr <= waddr;
        raddr <= raddr;
      end
    endcase
  end
end


endmodule
